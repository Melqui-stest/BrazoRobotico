-- Nombre: BRAZO_DEF - Structural
-- Con este c�digo se implementa el control conjunto de los servomotores y del motor paso a paso del brazo rob�tico dise�ado.
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
entity BRAZO_DEF is
  Port (
          clk : in std_logic;--Se�al de reloj de per�odo 10ns( mitad a 1 y mitad a 0)
          reset: in std_logic;--Reset del c�digo y se corresponde con el bot�n btnc de la FPGA.
  --------------------SERVOMOTOR
          --INPUTS
         --SW14 SW13 SW12 SW11 SW10-->Interruptores con los que se selecciona los servos correspondientes 
         -----------------------------a la articulaci�n en la que se quiera el movimiento.
          swselservos0 : in std_logic;    --SW10
          swselservos1 : in std_logic;    --SW11
          swselservos2 : in std_logic;    --SW12
          swselservos3 : in std_logic;    --SW13
          swselservos4 : in std_logic;    --SW14
          swgiroservos: in std_logic_vector(3 downto 0);--SW9 SW8 SW7 SW6-->Interruptores con los que se elige el angulo de giro del servo 
          ------swgiroservos----------Giro(�)
          --------0000------------------0---
          --------0001------------------18--
          --------0010------------------36--
          --------0011------------------54--
          --------0100------------------72--
          --------0101------------------90--
          --------0110------------------108--
          --------0111------------------126-
          --------1000------------------144-
          --------1001------------------162-
          --------1010------------------180-
          --OUTPUTS
          --JD5 JD4 JD3 JD2 JD1 JD0-->Puerto de salida por donde se obtiene la se�al de control de cada servo.
          ----------------------------Cada pin de salida JDi se corresponde  con la se�al de control de un servo diferente.
          JD0: out std_logic;--se�al de control servo 0
          JD1: out std_logic;--se�al de control servo 1
          JD2: out std_logic;--se�al de control servo 2
          JD3: out std_logic;--se�al de control servo 3
          JD4: out std_logic;--se�al de control servo 4
          JD5: out std_logic;--se�al de control servo 5
      
  --------------------STEPMOTOR
          --INPUTS
          swdir : in std_logic;--SW0-->Control de la direcci�n de giro.
          swenable: in std_logic;--SW5-->Interruptor enable--desactiva todo
          swoff: in std_logic;--SW4-->Activa o desactiva movimiento sin tocar el enable, por que si activas el enable deja de haber movimiento
          ----------------------------pero tambien fuerza desactiva movimiento pero mantiene fuerza.
          swgirostep: in std_logic_vector(2 downto 0);--SW3 SW2 SW1-->Interruptores con los que se ajusta el paso deseado(control del giro)
                          ---swgirostep    fincuenta     giro(�)
                          ---000    0              0
                          ---001    150.000      15
                          ---010    300.000      30
                          ---011    450.000      45
                          ---100    600.00       60
                          ---101    750.000      75
                          ---110    900.000      90
                          ---111    1.800.000    180
          --OUTPUTS
          enable: out std_logic;--JC1-->Se�al con la que se desactiva el motor
          dir: out std_logic; -- JC3-->Se�al con la que se establece el la direcci�n de giro del motor(0 en sentido horario y 1 en sentido antihorario)
          step : out std_logic --JC2-->Se�al peri�dica, con la que cada per�odo se consigue un giro del motor de un micropaso.
          -----------------------------En el caso en el que su valor sea cero, el giro del motor estar� desactivado. 
           );
end BRAZO_DEF;

architecture Structural of BRAZO_DEF is
component BRAZO_STEPMOTOR_DEF
 Port(
      clk : in std_logic;
      reset: in std_logic;-- ser� el reset(btnc)-btn0
      swdir : in std_logic;--control de la direcci�n--swt0
      swenable: in std_logic;--enable--desactiva todo
      swoff: in std_logic;--boton para activar o desactivar movimmiento sin tocar el enable, por que si activas el enable deja de haber movimiento pero tambien fuerza
     --desactiva movimiento pero mantiene fuerza
      swgirostep: in std_logic_vector(2 downto 0);--control del giro
      enable: out std_logic;--led0
      dir: out std_logic; -- 0 gira sentido horario y 1 sentido antihorario --led 4
      step : out std_logic -- se�al para cada micropaso--led5     
      );
 end component;
 
 component BRAZO_SERVOMOTOR_DEF
  Port(
       clk : in std_logic;
       reset: in std_logic;-- ser� el reset(btnc)-btn0
       swselservos0 : in std_logic;    --SW10
       swselservos1 : in std_logic;    --SW11
       swselservos2 : in std_logic;    --SW12
       swselservos3 : in std_logic;    --SW13
       swselservos4 : in std_logic;    --SW14
       swgiroservos: in std_logic_vector(3 downto 0);--ELECCION DE GIRO
       JD0: out std_logic;--se�al de control servo 0
       JD1: out std_logic;--se�al de control servo 1
       JD2: out std_logic;--se�al de control servo 2
       JD3: out std_logic;--se�al de control servo 3
       JD4: out std_logic;--se�al de control servo 4
       JD5: out std_logic--se�al de control servo 5
       );
  end component;
-----Servomotor
---- Inputs
--  signal clk : std_logic;
--  signal reset: std_logic;-- ser� el reset(btnc)
--  signal swselservos : std_logic_vector(5 downto 0);
--  signal  swgiroservos: std_logic_vector(3 downto 0);
--  --Outputs
--  signal JD: std_logic_vector( 5 downto 0);
----Stepmotor
----Inputps
----signal clk : std_logic;
----signal reset: std_logic;-- ser� el reset(btnc)
--signal swdir : std_logic;--control de la direcci�n(btnU)
--signal swenable: std_logic;--enable--desactiva todo
--signal swoff: std_logic;--enable--desactiva todo
--signal swgirostep:  std_logic_vector(2 downto 0);--control del giro
----Outputs
--signal  dir: std_logic; -- 0 gira sentido horario y 1 sentido antihorario --led 4
--signal step : std_logic; -- se�al para cada micropaso--led5
--signal enable: std_logic;--led0
begin
Portmap_stepmotor: BRAZO_STEPMOTOR_DEF
Port map (
            clk     =>  clk,
            reset   =>  reset,
            swdir  =>  swdir,
            swenable    =>  swenable,
            swoff    =>  swoff,
            swgirostep      =>  swgirostep,
            enable  =>  enable,
            dir     =>  dir,
            step    =>  step
          );
          
Portmap_servomotor: BRAZO_SERVOMOTOR_DEF
Port map (
            clk     =>  clk,
            reset   =>  reset,
            swselservos0     =>  swselservos0,
            swselservos1    =>  swselservos1,
            swselservos2     =>  swselservos2,
            swselservos3     =>  swselservos3,
            swselservos4     =>  swselservos4,
            swgiroservos     =>  swgiroservos,
            JD0      =>  JD0,
            JD1      =>  JD1,
            JD2      =>  JD2,
            JD3      =>  JD3,
            JD4      =>  JD4,
            JD5      =>  JD5
            
           );
end Structural;
